module fsm(input clk,input,rest,)